module main;
initial begin
    $display("Hello, World!\nThis is Verilog Programming Language.");
end
endmodule
